`include "sysarray16.v"
module sysarraytb16;

reg rst, clk;

reg [31:0] inp_west0, inp_west1, inp_west2, inp_west3, inp_west4, inp_west5, inp_west6, inp_west7, inp_west8, inp_west9, inp_west10, inp_west11, inp_west12, inp_west13, inp_west14, inp_west15, inp_north0, inp_north1, inp_north2, inp_north3, inp_north4, inp_north5, inp_north6, inp_north7, inp_north8, inp_north9, inp_north10, inp_north11, inp_north12, inp_north13, inp_north14, inp_north15;
wire okay;

sysarray16 uut16(inp_west0, inp_west1, inp_west2, inp_west3, inp_west4, inp_west5, inp_west6, inp_west7, inp_west8, inp_west9, inp_west10, inp_west11, inp_west12, inp_west13, inp_west14, inp_west15, inp_north0, inp_north1, inp_north2, inp_north3, inp_north4, inp_north5, inp_north6, inp_north7, inp_north8, inp_north9, inp_north10, inp_north11, inp_north12, inp_north13, inp_north14, inp_north15, 
		      clk, rst, fine);


initial begin
	#3  inp_west0 <= 32'd3;
	    inp_north0 <= 32'd12;
	#10 inp_west0 <= 32'd2;
	    inp_north0 <= 32'd8;
	#10 inp_west0 <= 32'd1;
	    inp_north0 <= 32'd4;
	#10 inp_west0 <= 32'd0;
	    inp_north0 <= 32'd0;
    #10 inp_west0 <= 32'd3;
	    inp_north0 <= 32'd12;
	#10 inp_west0 <= 32'd2;
	    inp_north0 <= 32'd8;
	#10 inp_west0 <= 32'd1;
	    inp_north0 <= 32'd4;
	#10 inp_west0 <= 32'd0;
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd3;
	    inp_north0 <= 32'd12;
	#10 inp_west0 <= 32'd2;
	    inp_north0 <= 32'd8;
	#10 inp_west0 <= 32'd1;
	    inp_north0 <= 32'd4;
	#10 inp_west0 <= 32'd0;
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd3;
	    inp_north0 <= 32'd12;
	#10 inp_west0 <= 32'd2;
	    inp_north0 <= 32'd8;
	#10 inp_west0 <= 32'd1;
	    inp_north0 <= 32'd4;
	#10 inp_west0 <= 32'd0;
	    inp_north0 <= 32'd0;
	#10 inp_west0 <= 32'd0;
	    inp_north0 <= 32'd0;
	#10 inp_west0 <= 32'd0;
	    inp_north0 <= 32'd0;
	#10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
        #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
        #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
        #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
        #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
         #10 inp_west0 <= 32'd0;	
	    inp_north0 <= 32'd0;
end

initial begin
	#3  inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
	#10 inp_west1 <= 32'd7;
	    inp_north1 <= 32'd13;
	#10 inp_west1 <= 32'd6;
	    inp_north1 <= 32'd9;
	#10 inp_west1 <= 32'd5;
	    inp_north1 <= 32'd5;
	#10 inp_west1 <= 32'd4;
	    inp_north1 <= 32'd1;
    #10 inp_west1 <= 32'd7;
	    inp_north1 <= 32'd13;
	#10 inp_west1 <= 32'd6;
	    inp_north1 <= 32'd9;
	#10 inp_west1 <= 32'd5;
	    inp_north1 <= 32'd5;
	#10 inp_west1 <= 32'd4;
	    inp_north1 <= 32'd1; 
    #10 inp_west1 <= 32'd7;
	    inp_north1 <= 32'd13;
	#10 inp_west1 <= 32'd6;
	    inp_north1 <= 32'd9;
	#10 inp_west1 <= 32'd5;
	    inp_north1 <= 32'd5;
	#10 inp_west1 <= 32'd4;
	    inp_north1 <= 32'd1;
        #10 inp_west1 <= 32'd7;
	    inp_north1 <= 32'd13;
	#10 inp_west1 <= 32'd6;
	    inp_north1 <= 32'd9;
	#10 inp_west1 <= 32'd5;
	    inp_north1 <= 32'd5;
	#10 inp_west1 <= 32'd4;
	    inp_north1 <= 32'd1;
    #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;           
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
	#10 inp_west1 <= 32'd0;
	    inp_north1 <= 32'd0;
	#10 inp_west1 <= 32'd0;	
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;	
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;	
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;	
	    inp_north1 <= 32'd0;
        #10 inp_west1 <= 32'd0;	
	    inp_north1 <= 32'd0;
end

initial begin
	#3  inp_west2 <= 32'd0;
	    inp_north2 <= 32'd0;
	#10 inp_west2 <= 32'd0;
	    inp_north2 <= 32'd0;
	#10 inp_west2 <= 32'd11;
	    inp_north2 <= 32'd14;
	#10 inp_west2 <= 32'd10;
	    inp_north2 <= 32'd10;
	#10 inp_west2 <= 32'd9;
	    inp_north2 <= 32'd6;
	#10 inp_west2 <= 32'd8;
	    inp_north2 <= 32'd2;
    #10 inp_west2 <= 32'd11;
	    inp_north2 <= 32'd14;
	#10 inp_west2 <= 32'd10;
	    inp_north2 <= 32'd10;
	#10 inp_west2 <= 32'd9;
	    inp_north2 <= 32'd6;
	#10 inp_west2 <= 32'd8;
	    inp_north2 <= 32'd2;
    #10 inp_west2 <= 32'd11;
	    inp_north2 <= 32'd14;
	#10 inp_west2 <= 32'd10;
	    inp_north2 <= 32'd10;
	#10 inp_west2 <= 32'd9;
	    inp_north2 <= 32'd6;
	#10 inp_west2 <= 32'd8;
	    inp_north2 <= 32'd2;
        #10 inp_west2 <= 32'd11;
	    inp_north2 <= 32'd14;
	#10 inp_west2 <= 32'd10;
	    inp_north2 <= 32'd10;
	#10 inp_west2 <= 32'd9;
	    inp_north2 <= 32'd6;
	#10 inp_west2 <= 32'd8;
	    inp_north2 <= 32'd2;        
	#10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
        #10 inp_west2 <= 32'd0;	
	    inp_north2 <= 32'd0;
end

initial begin
	#3  inp_west3 <= 32'd0;
	    inp_north3 <= 32'd0;
	#10 inp_west3 <= 32'd0;
	    inp_north3 <= 32'd0;
	#10 inp_west3 <= 32'd0;
	    inp_north3 <= 32'd0;
	#10 inp_west3 <= 32'd15;
	    inp_north3 <= 32'd15;
	#10 inp_west3 <= 32'd14;
	    inp_north3 <= 32'd11;
	#10 inp_west3 <= 32'd13;
	    inp_north3 <= 32'd7;
	#10 inp_west3 <= 32'd12;	
	    inp_north3 <= 32'd3;
    #10 inp_west3 <= 32'd15;
	    inp_north3 <= 32'd15;
	#10 inp_west3 <= 32'd14;
	    inp_north3 <= 32'd11;
	#10 inp_west3 <= 32'd13;
	    inp_north3 <= 32'd7;
	#10 inp_west3 <= 32'd12;	
	    inp_north3 <= 32'd3;
        #10 inp_west3 <= 32'd15;
	    inp_north3 <= 32'd15;
	#10 inp_west3 <= 32'd14;
	    inp_north3 <= 32'd11;
	#10 inp_west3 <= 32'd13;
	    inp_north3 <= 32'd7;
	#10 inp_west3 <= 32'd12;	
	    inp_north3 <= 32'd3;
        #10 inp_west3 <= 32'd15;
	    inp_north3 <= 32'd15;
	#10 inp_west3 <= 32'd14;
	    inp_north3 <= 32'd11;
	#10 inp_west3 <= 32'd13;
	    inp_north3 <= 32'd7;
	#10 inp_west3 <= 32'd12;	
	    inp_north3 <= 32'd3;   
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0; 
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0;
        #10 inp_west3 <= 32'd0;	
	    inp_north3 <= 32'd0; 
end

initial begin
	#3 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
        #10 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
        #10 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
        #10 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
    #10  inp_west4 <= 32'd3;
	    inp_north4 <= 32'd12;
	#10 inp_west4 <= 32'd2;
	    inp_north4 <= 32'd8;
	#10 inp_west4 <= 32'd1;
	    inp_north4 <= 32'd4;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
        #10  inp_west4 <= 32'd3;
	    inp_north4 <= 32'd12;
	#10 inp_west4 <= 32'd2;
	    inp_north4 <= 32'd8;
	#10 inp_west4 <= 32'd1;
	    inp_north4 <= 32'd4;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
    #10  inp_west4 <= 32'd3;
	    inp_north4 <= 32'd12;
	#10 inp_west4 <= 32'd2;
	    inp_north4 <= 32'd8;
	#10 inp_west4 <= 32'd1;
	    inp_north4 <= 32'd4;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
        #10  inp_west4 <= 32'd3;
	    inp_north4 <= 32'd12;
	#10 inp_west4 <= 32'd2;
	    inp_north4 <= 32'd8;
	#10 inp_west4 <= 32'd1;
	    inp_north4 <= 32'd4;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;    
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
    #10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
        #10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;	
	    inp_north4 <= 32'd0;
        #10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;
	#10 inp_west4 <= 32'd0;
	    inp_north4 <= 32'd0;    
end

initial begin
    #3 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
	#10 inp_west5 <= 32'd7;
	    inp_north5 <= 32'd13;
	#10 inp_west5 <= 32'd6;
	    inp_north5 <= 32'd9;
	#10 inp_west5 <= 32'd5;
	    inp_north5 <= 32'd5;
	#10 inp_west5 <= 32'd4;
	    inp_north5 <= 32'd1;
        #10 inp_west5 <= 32'd7;
	    inp_north5 <= 32'd13;
	#10 inp_west5 <= 32'd6;
	    inp_north5 <= 32'd9;
	#10 inp_west5 <= 32'd5;
	    inp_north5 <= 32'd5;
	#10 inp_west5 <= 32'd4;
	    inp_north5 <= 32'd1;
        #10 inp_west5 <= 32'd7;
	    inp_north5 <= 32'd13;
	#10 inp_west5 <= 32'd6;
	    inp_north5 <= 32'd9;
	#10 inp_west5 <= 32'd5;
	    inp_north5 <= 32'd5;
	#10 inp_west5 <= 32'd4;
	    inp_north5 <= 32'd1;
        #10 inp_west5 <= 32'd7;
	    inp_north5 <= 32'd13;
	#10 inp_west5 <= 32'd6;
	    inp_north5 <= 32'd9;
	#10 inp_west5 <= 32'd5;
	    inp_north5 <= 32'd5;
	#10 inp_west5 <= 32'd4;
	    inp_north5 <= 32'd1;
	#10 inp_west5 <= 32'd0;
	    inp_north5 <= 32'd0;
	#10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
        #10 inp_west5 <= 32'd0;	
	    inp_north5 <= 32'd0;
end

initial begin
	#3  inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
	#10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
	#10 inp_west6 <= 32'd11;
	    inp_north6 <= 32'd14;
	#10 inp_west6 <= 32'd10;
	    inp_north6 <= 32'd10;
	#10 inp_west6 <= 32'd9;
	    inp_north6 <= 32'd6;
	#10 inp_west6 <= 32'd8;
	    inp_north6 <= 32'd2;
        #10 inp_west6 <= 32'd11;
	    inp_north6 <= 32'd14;
	#10 inp_west6 <= 32'd10;
	    inp_north6 <= 32'd10;
	#10 inp_west6 <= 32'd9;
	    inp_north6 <= 32'd6;
	#10 inp_west6 <= 32'd8;
	    inp_north6 <= 32'd2;
           #10 inp_west6 <= 32'd11;
	    inp_north6 <= 32'd14;
	#10 inp_west6 <= 32'd10;
	    inp_north6 <= 32'd10;
	#10 inp_west6 <= 32'd9;
	    inp_north6 <= 32'd6;
	#10 inp_west6 <= 32'd8;
	    inp_north6 <= 32'd2;
           #10 inp_west6 <= 32'd11;
	    inp_north6 <= 32'd14;
	#10 inp_west6 <= 32'd10;
	    inp_north6 <= 32'd10;
	#10 inp_west6 <= 32'd9;
	    inp_north6 <= 32'd6;
	#10 inp_west6 <= 32'd8;
	    inp_north6 <= 32'd2;
	#10 inp_west6 <= 32'd0;	
	    inp_north6 <= 32'd0;
         #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
         #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
        #10 inp_west6 <= 32'd0;
	    inp_north6 <= 32'd0;
end

initial begin
	#3  inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
	#10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
	#10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
	#10 inp_west7 <= 32'd15;
	    inp_north7 <= 32'd15;
	#10 inp_west7 <= 32'd14;
	    inp_north7 <= 32'd11;
	#10 inp_west7 <= 32'd13;
	    inp_north7 <= 32'd7;
	#10 inp_west7 <= 32'd12;	
	    inp_north7 <= 32'd3;
        #10 inp_west7 <= 32'd15;
	    inp_north7 <= 32'd15;
	#10 inp_west7 <= 32'd14;
	    inp_north7 <= 32'd11;
	#10 inp_west7 <= 32'd13;
	    inp_north7 <= 32'd7;
	#10 inp_west7 <= 32'd12;	
	    inp_north7 <= 32'd3;
        #10 inp_west7 <= 32'd15;
	    inp_north7 <= 32'd15;
	#10 inp_west7 <= 32'd14;
	    inp_north7 <= 32'd11;
	#10 inp_west7 <= 32'd13;
	    inp_north7 <= 32'd7;
	#10 inp_west7 <= 32'd12;	
	    inp_north7 <= 32'd3;
        #10 inp_west7 <= 32'd15;
	    inp_north7 <= 32'd15;
	#10 inp_west7 <= 32'd14;
	    inp_north7 <= 32'd11;
	#10 inp_west7 <= 32'd13;
	    inp_north7 <= 32'd7;
	#10 inp_west7 <= 32'd12;	
	    inp_north7 <= 32'd3;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
        #10 inp_west7 <= 32'd0;
	    inp_north7 <= 32'd0;
end

initial begin
     #3 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;   
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0; 
         #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;   
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0; 
	#10  inp_west8 <= 32'd3;
	    inp_north8 <= 32'd12;
	#10 inp_west8 <= 32'd2;
	    inp_north8 <= 32'd8;
	#10 inp_west8 <= 32'd1;
	    inp_north8 <= 32'd4;
	#10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10  inp_west8 <= 32'd3;
	    inp_north8 <= 32'd12;
	#10 inp_west8 <= 32'd2;
	    inp_north8 <= 32'd8;
	#10 inp_west8 <= 32'd1;
	    inp_north8 <= 32'd4;
	#10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10  inp_west8 <= 32'd3;
	    inp_north8 <= 32'd12;
	#10 inp_west8 <= 32'd2;
	    inp_north8 <= 32'd8;
	#10 inp_west8 <= 32'd1;
	    inp_north8 <= 32'd4;
	#10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
    #10 inp_west8 <= 32'd3;
	    inp_north8 <= 32'd12;
	#10 inp_west8 <= 32'd2;
	    inp_north8 <= 32'd8;
	#10 inp_west8 <= 32'd1;
	    inp_north8 <= 32'd4;
	#10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
	#10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
	#10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
    #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;   
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0;
        #10 inp_west8 <= 32'd0;
	    inp_north8 <= 32'd0; 
end

initial begin
	#3  inp_west9 <= 32'd0;
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
	#10 inp_west9 <= 32'd7;
	    inp_north9 <= 32'd13;
	#10 inp_west9 <= 32'd6;
	    inp_north9 <= 32'd9;
	#10 inp_west9 <= 32'd5;
	    inp_north9 <= 32'd5;
	#10 inp_west9 <= 32'd4;
	    inp_north9 <= 32'd1;
        #10 inp_west9 <= 32'd7;
	    inp_north9 <= 32'd13;
	#10 inp_west9 <= 32'd6;
	    inp_north9 <= 32'd9;
	#10 inp_west9 <= 32'd5;
	    inp_north9 <= 32'd5;
	#10 inp_west9 <= 32'd4;
	    inp_north9 <= 32'd1;
        #10 inp_west9 <= 32'd7;
	    inp_north9 <= 32'd13;
	#10 inp_west9 <= 32'd6;
	    inp_north9 <= 32'd9;
	#10 inp_west9 <= 32'd5;
	    inp_north9 <= 32'd5;
	#10 inp_west9 <= 32'd4;
	    inp_north9 <= 32'd1;
    #10 inp_west9 <= 32'd7;
	    inp_north9 <= 32'd13;
	#10 inp_west9 <= 32'd6;
	    inp_north9 <= 32'd9;
	#10 inp_west9 <= 32'd5;
	    inp_north9 <= 32'd5;
	#10 inp_west9 <= 32'd4;
	    inp_north9 <= 32'd1;    
	#10 inp_west9 <= 32'd0;
	    inp_north9 <= 32'd0;
	#10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
        #10 inp_west9 <= 32'd0;	
	    inp_north9 <= 32'd0;
end

initial begin
	#3  inp_west10 <= 32'd0;
	    inp_north10 <= 32'd0;
         #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
         #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
	#10 inp_west10 <= 32'd0;
	    inp_north10 <= 32'd0;
	#10 inp_west10 <= 32'd11;
	    inp_north10 <= 32'd14;
	#10 inp_west10 <= 32'd10;
	    inp_north10 <= 32'd10;
	#10 inp_west10 <= 32'd9;
	    inp_north10 <= 32'd6;
	#10 inp_west10 <= 32'd8;
	    inp_north10 <= 32'd2;
        #10 inp_west10 <= 32'd11;
	    inp_north10 <= 32'd14;
	#10 inp_west10 <= 32'd10;
	    inp_north10 <= 32'd10;
	#10 inp_west10 <= 32'd9;
	    inp_north10 <= 32'd6;
	#10 inp_west10 <= 32'd8;
	    inp_north10 <= 32'd2;
        #10 inp_west10 <= 32'd11;
	    inp_north10 <= 32'd14;
	#10 inp_west10 <= 32'd10;
	    inp_north10 <= 32'd10;
	#10 inp_west10 <= 32'd9;
	    inp_north10 <= 32'd6;
	#10 inp_west10 <= 32'd8;
	    inp_north10 <= 32'd2;
    #10 inp_west10 <= 32'd11;
	    inp_north10 <= 32'd14;
	#10 inp_west10 <= 32'd10;
	    inp_north10 <= 32'd10;
	#10 inp_west10 <= 32'd9;
	    inp_north10 <= 32'd6;
	#10 inp_west10 <= 32'd8;
	    inp_north10 <= 32'd2;    
	#10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
        #10 inp_west10 <= 32'd0;	
	    inp_north10 <= 32'd0;
end

initial begin
	#3  inp_west11 <= 32'd0;
	    inp_north11 <= 32'd0;
         #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0; 
         #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0; 
	#10 inp_west11 <= 32'd0;
	    inp_north11 <= 32'd0;
	#10 inp_west11 <= 32'd0;
	    inp_north11 <= 32'd0;
	#10 inp_west11 <= 32'd15;
	    inp_north11 <= 32'd15;
	#10 inp_west11 <= 32'd14;
	    inp_north11 <= 32'd11;
	#10 inp_west11 <= 32'd13;
	    inp_north11 <= 32'd7;
	#10 inp_west11 <= 32'd12;	
	    inp_north11 <= 32'd3;
    #10 inp_west11 <= 32'd15;
	    inp_north11 <= 32'd15;
	#10 inp_west11 <= 32'd14;
	    inp_north11 <= 32'd11;
	#10 inp_west11 <= 32'd13;
	    inp_north11 <= 32'd7;
	#10 inp_west11 <= 32'd12;	
	    inp_north11 <= 32'd3;
        #10 inp_west11 <= 32'd15;
	    inp_north11 <= 32'd15;
	#10 inp_west11 <= 32'd14;
	    inp_north11 <= 32'd11;
	#10 inp_west11 <= 32'd13;
	    inp_north11 <= 32'd7;
	#10 inp_west11 <= 32'd12;	
	    inp_north11 <= 32'd3;  
        #10 inp_west11 <= 32'd15;
	    inp_north11 <= 32'd15;
	#10 inp_west11 <= 32'd14;
	    inp_north11 <= 32'd11;
	#10 inp_west11 <= 32'd13;
	    inp_north11 <= 32'd7;
	#10 inp_west11 <= 32'd12;	
	    inp_north11 <= 32'd3;     
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0;
        #10 inp_west11 <= 32'd0;	
	    inp_north11 <= 32'd0; 
end

initial begin
	#3 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
    #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
        #10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
    #10  inp_west12 <= 32'd3;
	    inp_north12 <= 32'd12;
	#10 inp_west12 <= 32'd2;
	    inp_north12 <= 32'd8;
	#10 inp_west12 <= 32'd1;
	    inp_north12 <= 32'd4;
	#10 inp_west12 <= 32'd0;
	    inp_north12 <= 32'd0;
       #10  inp_west12 <= 32'd3;
	    inp_north12 <= 32'd12;
	#10 inp_west12 <= 32'd2;
	    inp_north12 <= 32'd8;
	#10 inp_west12 <= 32'd1;
	    inp_north12 <= 32'd4;
	#10 inp_west12 <= 32'd0;
	    inp_north12 <= 32'd0;
        #10  inp_west12 <= 32'd3;
	    inp_north12 <= 32'd12;
	#10 inp_west12 <= 32'd2;
	    inp_north12 <= 32'd8;
	#10 inp_west12 <= 32'd1;
	    inp_north12 <= 32'd4;
	#10 inp_west12 <= 32'd0;
	    inp_north12 <= 32'd0;
        #10  inp_west12 <= 32'd3;
	    inp_north12 <= 32'd12;
	#10 inp_west12 <= 32'd2;
	    inp_north12 <= 32'd8;
	#10 inp_west12 <= 32'd1;
	    inp_north12 <= 32'd4;
	#10 inp_west12 <= 32'd0;
	    inp_north12 <= 32'd0;
	#10 inp_west12 <= 32'd0;
	    inp_north12 <= 32'd0;
	#10 inp_west12 <= 32'd0;
	    inp_north12 <= 32'd0;
	#10 inp_west12 <= 32'd0;	
	    inp_north12 <= 32'd0;
end

initial begin
    #3 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
       #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
        #10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
	#10 inp_west13 <= 32'd7;
	    inp_north13 <= 32'd13;
	#10 inp_west13 <= 32'd6;
	    inp_north13 <= 32'd9;
	#10 inp_west13 <= 32'd5;
	    inp_north13 <= 32'd5;
	#10 inp_west13 <= 32'd4;
	    inp_north13 <= 32'd1;
#10 inp_west13 <= 32'd7;
	    inp_north13 <= 32'd13;
	#10 inp_west13 <= 32'd6;
	    inp_north13 <= 32'd9;
	#10 inp_west13 <= 32'd5;
	    inp_north13 <= 32'd5;
	#10 inp_west13 <= 32'd4;
	    inp_north13 <= 32'd1;
        #10 inp_west13 <= 32'd7;
	    inp_north13 <= 32'd13;
	#10 inp_west13 <= 32'd6;
	    inp_north13 <= 32'd9;
	#10 inp_west13 <= 32'd5;
	    inp_north13 <= 32'd5;
	#10 inp_west13 <= 32'd4;
	    inp_north13 <= 32'd1;
        #10 inp_west13 <= 32'd7;
	    inp_north13 <= 32'd13;
	#10 inp_west13 <= 32'd6;
	    inp_north13 <= 32'd9;
	#10 inp_west13 <= 32'd5;
	    inp_north13 <= 32'd5;
	#10 inp_west13 <= 32'd4;
	    inp_north13 <= 32'd1;
	#10 inp_west13 <= 32'd0;
	    inp_north13 <= 32'd0;
	#10 inp_west13 <= 32'd0;	
	    inp_north13 <= 32'd0;
end

initial begin
	#3  inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
       #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
	#10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
         #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
	#10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
         #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
        #10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
	#10 inp_west14 <= 32'd0;
	    inp_north14 <= 32'd0;
	#10 inp_west14 <= 32'd11;
	    inp_north14 <= 32'd14;
	#10 inp_west14 <= 32'd10;
	    inp_north14 <= 32'd10;
	#10 inp_west14 <= 32'd9;
	    inp_north14 <= 32'd6;
	#10 inp_west14 <= 32'd8;
	    inp_north14 <= 32'd2;
        #10 inp_west14 <= 32'd11;
	    inp_north14 <= 32'd14;
	#10 inp_west14 <= 32'd10;
	    inp_north14 <= 32'd10;
	#10 inp_west14 <= 32'd9;
	    inp_north14 <= 32'd6;
	#10 inp_west14 <= 32'd8;
	    inp_north14 <= 32'd2;
        #10 inp_west14 <= 32'd11;
	    inp_north14 <= 32'd14;
	#10 inp_west14 <= 32'd10;
	    inp_north14 <= 32'd10;
	#10 inp_west14 <= 32'd9;
	    inp_north14 <= 32'd6;
	#10 inp_west14 <= 32'd8;
	    inp_north14 <= 32'd2;
        #10 inp_west14 <= 32'd11;
	    inp_north14 <= 32'd14;
	#10 inp_west14 <= 32'd10;
	    inp_north14 <= 32'd10;
	#10 inp_west14 <= 32'd9;
	    inp_north14 <= 32'd6;
	#10 inp_west14 <= 32'd8;
	    inp_north14 <= 32'd2;
	#10 inp_west14 <= 32'd0;	
	    inp_north14 <= 32'd0;
end

initial begin
	#3  inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
	#10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
        #10 inp_west15 <= 32'd0;
	    inp_north15 <= 32'd0;
	#10 inp_west15 <= 32'd15;
	    inp_north15 <= 32'd15;
	#10 inp_west15 <= 32'd14;
	    inp_north15 <= 32'd11;
	#10 inp_west15 <= 32'd13;
	    inp_north15 <= 32'd7;
	#10 inp_west15 <= 32'd12;	
	    inp_north15 <= 32'd3;
        #10 inp_west15 <= 32'd15;
	    inp_north15 <= 32'd15;
	#10 inp_west15 <= 32'd14;
	    inp_north15 <= 32'd11;
	#10 inp_west15 <= 32'd13;
	    inp_north15 <= 32'd7;
	#10 inp_west15 <= 32'd12;	
	    inp_north15 <= 32'd3;
        #10 inp_west15 <= 32'd15;
	    inp_north15 <= 32'd15;
	#10 inp_west15 <= 32'd14;
	    inp_north15 <= 32'd11;
	#10 inp_west15 <= 32'd13;
	    inp_north15 <= 32'd7;
	#10 inp_west15 <= 32'd12;	
	    inp_north15 <= 32'd3;
        #10 inp_west15 <= 32'd15;
	    inp_north15 <= 32'd15;
	#10 inp_west15 <= 32'd14;
	    inp_north15 <= 32'd11;
	#10 inp_west15 <= 32'd13;
	    inp_north15 <= 32'd7;
	#10 inp_west15 <= 32'd12;	
	    inp_north15 <= 32'd3;
end

initial 
begin
$monitor ($time,"East0=%b, East1=%b, East2=%b, East3=%b, East4=%b, East5=%b, East6=%b, East7=%b, East8=%b, East9=%b, East10=%b, East11=%b, East12=%b, East13=%b, East14=%b, East15=%b", uut16.reseast0, uut16.reseast1, uut16.reseast2, uut16.reseast3, uut16.reseast4, uut16.reseast5, uut16.reseast6, uut16.reseast7, uut16.reseast8, uut16.reseast9, uut16.reseast10, uut16.reseast11, uut16.reseast12, uut16.reseast13, uut16.reseast14, uut16.reseast15);
end

initial begin
rst <= 1;
clk <= 0;
#3
rst <= 0;
end

initial begin
	repeat(100)
		#5 clk <= ~clk;
end




initial begin
	$dumpfile("wave16.vcd");
	$dumpvars(0, sysarraytb16);
end



endmodule